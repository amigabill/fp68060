-- This is the top-level of the fp68060 design, instantiating
-- all top IP blocks, connecting things to external FPGA pins



